/*
TESTASE 2
*/